package Constants;
    localparam int unsigned BYTE           = 8;
    localparam int unsigned WIDTH          = 32;
    localparam int unsigned REG_ADDR_WIDTH = 5;
    localparam int unsigned REG_COUNT      = 32;
    localparam int unsigned ROM_SIZE       = 2 * 1024;
    localparam int unsigned RAM_SIZE       = 128;
    localparam int unsigned TARGET_WIDTH   = 26;
    localparam int unsigned SHAMT_WIDTH    = 5;
    localparam int unsigned IMM_WIDTH      = 16;
endpackage