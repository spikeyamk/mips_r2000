// Register Arithmetic Operations:
localparam Mask ADD    = 32'b000000???????????????00000100000;
localparam Mask ADDU   = 32'b000000???????????????00000100001;
localparam Mask SUB    = 32'b000000???????????????00000100010;
localparam Mask SUBU   = 32'b000000???????????????00000100011;
// Register Logic Operations:
localparam Mask AND    = 32'b000000???????????????00000100100;
localparam Mask OR     = 32'b000000???????????????00000100101;
localparam Mask XOR    = 32'b000000???????????????00000100110;
localparam Mask NOR    = 32'b000000???????????????00000100111;
// Register Shift Operations:
localparam Mask SLL    = 32'b00000000000???????????????000000;
localparam Mask SRL    = 32'b00000000000???????????????000010;
localparam Mask SRA    = 32'b00000000000???????????????000011;
localparam Mask SLLV   = 32'b000000???????????????00000000100;
localparam Mask SRLV   = 32'b000000???????????????00000000110;
localparam Mask SRAV   = 32'b000000???????????????00000000111;
// Register Comparison Operations:
localparam Mask SLT    = 32'b000000???????????????00000101010;
localparam Mask SLTU   = 32'b000000???????????????00000101011;
// Immediate Arithmetic Operations:
localparam Mask ADDI   = 32'b001000??????????????????????????;
localparam Mask ADDIU  = 32'b001001??????????????????????????;
// Immediate Logic Operations:
localparam Mask ANDI   = 32'b001100??????????????????????????;
localparam Mask ORI    = 32'b001101??????????????????????????;
localparam Mask XORI   = 32'b001110??????????????????????????;
// Immediate Comparison Operations:
localparam Mask SLTI   = 32'b001010??????????????????????????;
localparam Mask SLTIU  = 32'b001011??????????????????????????;
// Load and Store Operations:
localparam Mask LUI    = 32'b00111100000?????????????????????;
localparam Mask LB     = 32'b100000??????????????????????????;
localparam Mask LBU    = 32'b100100??????????????????????????;
localparam Mask LH     = 32'b100001??????????????????????????;
localparam Mask LHU    = 32'b100101??????????????????????????;
localparam Mask LW     = 32'b100011??????????????????????????;
localparam Mask LD     = 32'b110111??????????????????????????;
localparam Mask SB     = 32'b101000??????????????????????????;
localparam Mask SH     = 32'b101001??????????????????????????;
localparam Mask SW     = 32'b101011??????????????????????????;
localparam Mask SD     = 32'b111111??????????????????????????;
// Branch Operations:
localparam Mask BEQ    = 32'b000100??????????????????????????;
localparam Mask BNE    = 32'b000101??????????????????????????;
localparam Mask BLTZ   = 32'b000001?????00000????????????????;
localparam Mask BGEZ   = 32'b000001?????00001????????????????;
localparam Mask BLTZAL = 32'b000001?????10000????????????????;
localparam Mask BGEZAL = 32'b000001?????10001????????????????;
localparam Mask BLEZ   = 32'b000110?????00000????????????????;
localparam Mask BGTZ   = 32'b000111?????00000????????????????;
// Jump Operations:
localparam Mask J      = 32'b000010??????????????????????????;
localparam Mask JAL    = 32'b000011??????????????????????????;
localparam Mask JR     = 32'b000000?????000000000000000001000;
localparam Mask JALR   = 32'b000000?????00000?????00000001001;